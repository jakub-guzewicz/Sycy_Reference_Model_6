module hulkFinder(
	input clk,
	input ena,
	input rst,
	input mode,
	input [63:0] cipher,
	output [127:0] cipherKey
	
	);
	
	//REG/WIRE
	wire	[29:0] lfsr;
	wire	[7:0] char0;
	wire	[7:0] char1;
	wire	[7:0] char2;
	wire	[7:0] char3;
	wire	[7:0] char4;
	wire	[7:0] char5;
	wire	[127:0] key;
	wire	[63:0] decrypted;
	reg	[79:0] firstKeyPart;
	
	always@(mode)
	begin
		if(mode==1'b0)
			firstKeyPart = 80'h48756c6b206973207468;
		else
			firstKeyPart = 80'h48554c4b204953205448;
	end
	
	assign key = {firstKeyPart,char5,char4,char3,char2,char1,char0};
	
	random_generator gen0(
		.rst	(rst),
		.clk	(clk),
		.ena	(ena),
		.lfsr_next(lfsr)
		
	);
	
	fiveBitToAsciiDecoder dec0(
		.data(lfsr[4:0]),
		.mode(mode),
		.char(char0)
	);
	
	fiveBitToAsciiDecoder dec1(
		.data(lfsr[9:5]),
		.mode(mode),
		.char(char1)
	);
	
	fiveBitToAsciiDecoder dec2(
		.data(lfsr[14:10]),
		.mode(mode),
		.char(char2)
	);
	
	fiveBitToAsciiDecoder dec3(
		.data(lfsr[19:15]),
		.mode(mode),
		.char(char3)
	);
	
	fiveBitToAsciiDecoder dec4(
		.data(lfsr[24:20]),
		.mode(mode),
		.char(char4)
	);
	
	fiveBitToAsciiDecoder dec5(
		.data(lfsr[29:25]),
		.mode(mode),
		.char(char5)
	);
	
// First version
/*	teaDecryptor tea0(
		.cipher(cipher),
		.key(key),
		.data(decrypted)
	);
*/
	pdfCheckerFsm fsm0(
		.rst(rst),
		.clk(clk),
		.ena(ena),
		.givenKey(key),
		.data(decrypted),
		.foundKey(cipherKey)		
	);
//Second version D:
//	with wires

	wire [63:0] teaWire01;
	wire [63:0] teaWire12;
	wire [63:0] teaWire23;
	wire [63:0] teaWire34;
	wire [63:0] teaWire45;
	wire [63:0] teaWire56;
	wire [63:0] teaWire67;
	wire [63:0] teaWire78;
	wire [63:0] teaWire89;
	wire [63:0] teaWire910;
	wire [63:0] teaWire1011;
	wire [63:0] teaWire1112;
	wire [63:0] teaWire1213;
	wire [63:0] teaWire1314;
	wire [63:0] teaWire1415;
	wire [63:0] teaWire1516;
	wire [63:0] teaWire1617;
	wire [63:0] teaWire1718;
	wire [63:0] teaWire1819;
	wire [63:0] teaWire1920;
	wire [63:0] teaWire2021;
	wire [63:0] teaWire2122;
	wire [63:0] teaWire2223;
	wire [63:0] teaWire2324;
	wire [63:0] teaWire2425;
	wire [63:0] teaWire2526;
	wire [63:0] teaWire2627;
	wire [63:0] teaWire2728;
	wire [63:0] teaWire2829;
	wire [63:0] teaWire2930;
	wire [63:0] teaWire3031;
	wire [63:0] teaWire3132;

	
	singleTeaBlock tea0(
		.key(key),
		.clk(clk),
		.inData(cipher),
		.sum(32'hc6ef3720),
		.outData(teaWire01)
	);

	singleTeaBlock tea1(
		.key(key),
		.clk(clk),
		.inData(teaWire01),
		.sum(32'h28b7bd67),
		.outData(teaWire12)
	);

	singleTeaBlock tea2(
		.key(key),
		.clk(clk),
		.inData(teaWire12),
		.sum(32'h8a8043ae),
		.outData(teaWire23)
	);

	singleTeaBlock tea3(
		.key(key),
		.clk(clk),
		.inData(teaWire23),
		.sum(32'hec48c9f5),
		.outData(teaWire34)
	);

	singleTeaBlock tea4(
		.key(key),
		.clk(clk),
		.inData(teaWire34),
		.sum(32'h4e11503c),
		.outData(teaWire45)
	);

	singleTeaBlock tea5(
		.key(key),
		.clk(clk),
		.inData(teaWire45),
		.sum(32'hafd9d683),
		.outData(teaWire56)
	);

	singleTeaBlock tea6(
		.key(key),
		.clk(clk),
		.inData(teaWire56),
		.sum(32'h11a25cca),
		.outData(teaWire67)
	);

	singleTeaBlock tea7(
		.key(key),
		.clk(clk),
		.inData(teaWire67),
		.sum(32'h736ae311),
		.outData(teaWire78)
	);

	singleTeaBlock tea8(
		.key(key),
		.clk(clk),
		.inData(teaWire78),
		.sum(32'hd5336958),
		.outData(teaWire89)
	);

	singleTeaBlock tea9(
		.key(key),
		.clk(clk),
		.inData(teaWire89),
		.sum(32'h36fbef9f),
		.outData(teaWire910)
	);

	singleTeaBlock tea10(
		.key(key),
		.clk(clk),
		.inData(teaWire910),
		.sum(32'h98c475e6),
		.outData(teaWire1011)
	);

	singleTeaBlock tea11(
		.key(key),
		.clk(clk),
		.inData(teaWire1011),
		.sum(32'hfa8cfc2d),
		.outData(teaWire1112)
	);

	singleTeaBlock tea12(
		.key(key),
		.clk(clk),
		.inData(teaWire1112),
		.sum(32'h5c558274),
		.outData(teaWire1213)
	);

	singleTeaBlock tea13(
		.key(key),
		.clk(clk),
		.inData(teaWire1213),
		.sum(32'hbe1e08bb),
		.outData(teaWire1314)
	);

	singleTeaBlock tea14(
		.key(key),
		.clk(clk),
		.inData(teaWire1314),
		.sum(32'h1fe68f02),
		.outData(teaWire1415)
	);

	singleTeaBlock tea15(
		.key(key),
		.clk(clk),
		.inData(teaWire1415),
		.sum(32'h81af1549),
		.outData(teaWire1516)
	);

	singleTeaBlock tea16(
		.key(key),
		.clk(clk),
		.inData(teaWire1516),
		.sum(32'he3779b90),
		.outData(teaWire1617)
	);

	singleTeaBlock tea17(
		.key(key),
		.clk(clk),
		.inData(teaWire1617),
		.sum(32'h454021d7),
		.outData(teaWire1718)
	);

	singleTeaBlock tea18(
		.key(key),
		.clk(clk),
		.inData(teaWire1718),
		.sum(32'ha708a81e),
		.outData(teaWire1819)
	);

	singleTeaBlock tea19(
		.key(key),
		.clk(clk),
		.inData(teaWire1819),
		.sum(32'h8d12e65),
		.outData(teaWire1920)
	);

	singleTeaBlock tea20(
		.key(key),
		.clk(clk),
		.inData(teaWire1920),
		.sum(32'h6a99b4ac),
		.outData(teaWire2021)
	);

	singleTeaBlock tea21(
		.key(key),
		.clk(clk),
		.inData(teaWire2021),
		.sum(32'hcc623af3),
		.outData(teaWire2122)
	);

	singleTeaBlock tea22(
		.key(key),
		.clk(clk),
		.inData(teaWire2122),
		.sum(32'h2e2ac13a),
		.outData(teaWire2223)
	);

	singleTeaBlock tea23(
		.key(key),
		.clk(clk),
		.inData(teaWire2223),
		.sum(32'h8ff34781),
		.outData(teaWire2324)
	);

	singleTeaBlock tea24(
		.key(key),
		.clk(clk),
		.inData(teaWire2324),
		.sum(32'hf1bbcdc8),
		.outData(teaWire2425)
	);

	singleTeaBlock tea25(
		.key(key),
		.clk(clk),
		.inData(teaWire2425),
		.sum(32'h5384540f),
		.outData(teaWire2526)
	);

	singleTeaBlock tea26(
		.key(key),
		.clk(clk),
		.inData(teaWire2526),
		.sum(32'hb54cda56),
		.outData(teaWire2627)
	);

	singleTeaBlock tea27(
		.key(key),
		.clk(clk),
		.inData(teaWire2627),
		.sum(32'h1715609d),
		.outData(teaWire2728)
	);

	singleTeaBlock tea28(
		.key(key),
		.clk(clk),
		.inData(teaWire2728),
		.sum(32'h78dde6e4),
		.outData(teaWire2829)
	);

	singleTeaBlock tea29(
		.clk(clk),
		.key(key),
		.inData(teaWire2829),
		.sum(32'hdaa66d2b),
		.outData(teaWire2930)
	);

	singleTeaBlock tea30(
		.clk(clk),
		.key(key),
		.inData(teaWire2930),
		.sum(32'h3c6ef372),
		.outData(teaWire3031)
	);

	singleTeaBlock tea31(
		.clk(clk),
		.key(key),
		.inData(teaWire3031),
		.sum(32'h9e3779b9),
		.outData(decrypted)
	);

endmodule